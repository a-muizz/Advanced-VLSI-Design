module FIR_Filter_L3_Top 
#(
    parameter DATA_IN_WIDTH  = 16,
    parameter DATA_OUT_WIDTH = 64,
    parameter TAP_WIDTH      = 24,
    parameter TAP_COUNT      = 36
)
(
    input wire                               clk,
    input wire                               reset_n,
    input wire   signed [DATA_IN_WIDTH-1:0]  data_in_1,
	 input wire   signed [DATA_IN_WIDTH-1:0]  data_in_2,
	 input wire   signed [DATA_IN_WIDTH-1:0]  data_in_3,
    output reg   signed [DATA_OUT_WIDTH-1:0] data_out_1,
	 output reg   signed [DATA_OUT_WIDTH-1:0] data_out_2,
	 output reg   signed [DATA_OUT_WIDTH-1:0] data_out_3
);

//input side of diagram
reg [DATA_IN_WIDTH-1:0] data_input_H0H1, data_input_H1H2, data_input_H0H1H2;
assign data_input_H0H1 = data_in_1 + data_in_2;
assign data_input_H1H2 = data_in_2 + data_in_3;
assign data_input_H0H1H2 = data_input_H0H1 + data_in_3;


//Data out for sub parallel filters
reg [DATA_OUT_WIDTH-1:0] dataOut_H0, dataOut_H1, dataOut_H2, dataOut_H0H1, dataOut_H1H2, dataOut_H0H1H2;


// Tap coefficients (Paste generated tap values here)
localparam signed [TAP_WIDTH-1:0] H0_taps [0:TAP_COUNT-1] = '{24'b000000000000010010001100, 24'b000000000010010111000001, 24'b111111111101100101100110, 24'b111111011000100111111010, 24'b111110011110111101100101, 24'b111110100100110100101100, 24'b000000000010110111000100, 24'b000000110011110111101110, 24'b111111110100000111100101, 24'b111111011001000100000100, 24'b000000011011101010000010, 24'b000000010111000001111110, 24'b111111010011100100000110, 24'b000000000100101011001010, 24'b000000110111100010100001, 24'b111111000110101010111101, 24'b111111010000000110001001, 24'b000100000101011001111110, 24'b000110011101101101110000, 24'b000010010000110000001000, 24'b111110100110101110000101, 24'b111111110100110010001000, 24'b000000111000010001110110, 24'b111111100110011011101100, 24'b111111100011100010001000, 24'b000000100111011110101001, 24'b000000000100010000000111, 24'b111111010100001001011011, 24'b000000001111001000011100, 24'b000000110001110001100011, 24'b111111011111111001001101, 24'b111110010110110010010110, 24'b111110110000000100110101, 24'b111111101001100000111101, 24'b000000000001011100010010, 24'b000000000001100011011110};

localparam signed [TAP_WIDTH-1:0] H1_taps [0:TAP_COUNT-1] = '{24'b000000000000110001111111, 24'b000000000010101000100000, 24'b111111110101110111110011, 24'b111111000100100100001011, 24'b111110010101011000011000, 24'b111110111110011111001000, 24'b000000100000001111100100, 24'b000000100110110110110100, 24'b111111011110001100000000, 24'b111111101011001010010100, 24'b000000101001000100110101, 24'b111111111101010010110111, 24'b111111010100001100000001, 24'b000000100100000111001000, 24'b000000011111000011010110, 24'b111110100110111101110100, 24'b000000100010010100111110, 24'b000101100110100100101110, 24'b000101100110100100101110, 24'b000000100010010100111110, 24'b111110100110111101110100, 24'b000000011111000011010110, 24'b000000100100000111001000, 24'b111111010100001100000001, 24'b111111111101010010110111, 24'b000000101001000100110101, 24'b111111101011001010010100, 24'b111111011110001100000000, 24'b000000100110110110110100, 24'b000000100000001111100100, 24'b111110111110011111001000, 24'b111110010101011000011000, 24'b111111000100100100001011, 24'b111111110101110111110011, 24'b000000000010101000100000, 24'b000000000000110001111111};

localparam signed [TAP_WIDTH-1:0] H2_taps [0:TAP_COUNT-1] = '{24'b000000000001100011011110, 24'b000000000001011100010010, 24'b111111101001100000111101, 24'b111110110000000100110101, 24'b111110010110110010010110, 24'b111111011111111001001101, 24'b000000110001110001100011, 24'b000000001111001000011100, 24'b111111010100001001011011, 24'b000000000100010000000111, 24'b000000100111011110101001, 24'b111111100011100010001000, 24'b111111100110011011101100, 24'b000000111000010001110110, 24'b111111110100110010001000, 24'b111110100110101110000101, 24'b000010010000110000001000, 24'b000110011101101101110000, 24'b000100000101011001111110, 24'b111111010000000110001001, 24'b111111000110101010111101, 24'b000000110111100010100001, 24'b000000000100101011001010, 24'b111111010011100100000110, 24'b000000010111000001111110, 24'b000000011011101010000010, 24'b111111011001000100000100, 24'b111111110100000111100101, 24'b000000110011110111101110, 24'b000000000010110111000100, 24'b111110100100110100101100, 24'b111110011110111101100101, 24'b111111011000100111111010, 24'b111111111101100101100110, 24'b000000000010010111000001, 24'b000000000000010010001100};

localparam signed [TAP_WIDTH-1:0] H0_H1_taps [0:TAP_COUNT-1] = '{24'b000000000001000100001011, 24'b000000000100111111100001, 24'b111111110011011101011001, 24'b111110011101001100000101, 24'b111100110100010101111101, 24'b111101100011010011110100, 24'b000000100011000110101000, 24'b000001011010101110100010, 24'b111111010010010011100101, 24'b111111000100001110011000, 24'b000001000100101110110111, 24'b000000010100010100110101, 24'b111110100111110000000111, 24'b000000101000110010010010, 24'b000001010110100101110111, 24'b111101101101101000110001, 24'b111111110010011011000111, 24'b001001101011111110101100, 24'b001100000100010010011110, 24'b000010110011000101000110, 24'b111101001101101011111001, 24'b000000010011110101011110, 24'b000001011100011000111110, 24'b111110111010100111101101, 24'b111111100000110100111111, 24'b000001010000100011011110, 24'b111111101111011010011011, 24'b111110110010010101011011, 24'b000000110101111111010000, 24'b000001010010000001000111, 24'b111110011110011000010101, 24'b111100101100001010101110, 24'b111101110100101001000000, 24'b111111011111011000110000, 24'b000000000100000100110010, 24'b000000000010010101011101};

localparam signed [TAP_WIDTH-1:0] H1_H2_taps [0:TAP_COUNT-1] = '{24'b000000000010010101011101, 24'b000000000100000100110010, 24'b111111011111011000110000, 24'b111101110100101001000000, 24'b111100101100001010101110, 24'b111110011110011000010101, 24'b000001010010000001000111, 24'b000000110101111111010000, 24'b111110110010010101011011, 24'b111111101111011010011011, 24'b000001010000100011011110, 24'b111111100000110100111111, 24'b111110111010100111101101, 24'b000001011100011000111110, 24'b000000010011110101011110, 24'b111101001101101011111001, 24'b000010110011000101000110, 24'b001100000100010010011110, 24'b001001101011111110101100, 24'b111111110010011011000111, 24'b111101101101101000110001, 24'b000001010110100101110111, 24'b000000101000110010010010, 24'b111110100111110000000111, 24'b000000010100010100110101, 24'b000001000100101110110111, 24'b111111000100001110011000, 24'b111111010010010011100101, 24'b000001011010101110100010, 24'b000000100011000110101000, 24'b111101100011010011110100, 24'b111100110100010101111101, 24'b111110011101001100000101, 24'b111111110011011101011001, 24'b000000000100111111100001, 24'b000000000001000100001011};

localparam signed [TAP_WIDTH-1:0] H0_H1_H2_taps [0:TAP_COUNT-1] = '{24'b000000000010100111101001, 24'b000000000110011011110011, 24'b111111011100111110010110, 24'b111101001101010000111010, 24'b111011001011001000010011, 24'b111101000011001101000001, 24'b000001010100111000001011, 24'b000001101001110110111110, 24'b111110100110011101000000, 24'b111111001000011110011111, 24'b000001101100001101100000, 24'b111111110111110110111101, 24'b111110001110001011110011, 24'b000001100001000100001000, 24'b000001001011010111111111, 24'b111100010100010110110110, 24'b000010000011001011001111, 24'b010000001001101100011100, 24'b010000001001101100011100, 24'b000010000011001011001111, 24'b111100010100010110110110, 24'b000001001011010111111111, 24'b000001100001000100001000, 24'b111110001110001011110011, 24'b111111110111110110111101, 24'b000001101100001101100000, 24'b111111001000011110011111, 24'b111110100110011101000000, 24'b000001101001110110111110, 24'b000001010100111000001011, 24'b111101000011001101000001, 24'b111011001011001000010011, 24'b111101001101010000111010, 24'b111111011100111110010110, 24'b000000000110011011110011, 24'b000000000010100111101001};





fir_pipeline #( .TAPS(H0_taps) ) H0(clk, reset_n, data_in_1, dataOut_H0);
fir_pipeline #( .TAPS(H1_taps) ) H1(clk, reset_n, data_in_2, dataOut_H1);
fir_pipeline #( .TAPS(H2_taps) ) H2(clk, reset_n, data_in_3, dataOut_H2);
fir_pipeline #( .TAPS(H0_H1_taps) ) H0_H1(clk, reset_n, data_input_H0H1, dataOut_H0H1);
fir_pipeline #( .TAPS(H1_H2_taps) ) H1_H2(clk, reset_n, data_input_H1H2, dataOut_H1H2);
fir_pipeline #( .TAPS(H0_H1_H2_taps) ) H0_H1_H2(clk, reset_n, data_input_H0H1H2, dataOut_H0H1H2);


//output side of diagram:
reg signed [DATA_OUT_WIDTH-1:0] H2delay;
reg signed [DATA_OUT_WIDTH-1:0] H1_H1H2delay;
integer i;
//-----------------------------------------------------------
// Delay Line (for H1)
//-----------------------------------------------------------
always @(posedge clk or negedge reset_n) begin
    if (!reset_n) begin
       
            H2delay <= 0;
				H1_H1H2delay <= 0;
		
    end else begin
        // Shift the delay line: new sample enters at delay[0]
        
        H2delay <= dataOut_H2;
		  H1_H1H2delay <= dataOut_H1H2 - dataOut_H1;
    end
end


assign data_out_1 = dataOut_H0 - H2delay + H1_H1H2delay;
assign data_out_2 = dataOut_H0H1 - dataOut_H1 - (dataOut_H0 - H2delay);
assign data_out_3 = dataOut_H0H1H2 - (dataOut_H0H1 - dataOut_H1) - (dataOut_H1H2 - dataOut_H1);

endmodule