module fir_pipeline 
#(
    parameter DATA_IN_WIDTH  = 16,
    parameter DATA_OUT_WIDTH = 64,
    parameter TAP_WIDTH      = 24,
    parameter TAP_COUNT      = 108
)
(
    input wire                               clk,
    input wire                               reset_n,
    input wire   signed [DATA_IN_WIDTH-1:0]  data_in,
    output reg   signed [DATA_OUT_WIDTH-1:0] data_out
);

//-----------------------------------------------------------
// Internal registers and arrays
//-----------------------------------------------------------

// Delay line for input samples
reg signed [DATA_IN_WIDTH-1:0] delay [0:TAP_COUNT-1];

// Coefficient values for each tap
reg signed [TAP_WIDTH-1:0]  taps [0:TAP_COUNT-1] = '{24'b000000000000010010001100, 24'b000000000000110001111111, 24'b000000000001100011011110, 24'b000000000010010111000001, 24'b000000000010101000100000, 24'b000000000001011100010010, 24'b111111111101100101100110, 24'b111111110101110111110011, 24'b111111101001100000111101, 24'b111111011000100111111010, 24'b111111000100100100001011, 24'b111110110000000100110101, 24'b111110011110111101100101, 24'b111110010101011000011000, 24'b111110010110110010010110, 24'b111110100100110100101100, 24'b111110111110011111001000, 24'b111111011111111001001101, 24'b000000000010110111000100, 24'b000000100000001111100100, 24'b000000110001110001100011, 24'b000000110011110111101110, 24'b000000100110110110110100, 24'b000000001111001000011100, 24'b111111110100000111100101, 24'b111111011110001100000000, 24'b111111010100001001011011, 24'b111111011001000100000100, 24'b111111101011001010010100, 24'b000000000100010000000111, 24'b000000011011101010000010, 24'b000000101001000100110101, 24'b000000100111011110101001, 24'b000000010111000001111110, 24'b111111111101010010110111, 24'b111111100011100010001000, 24'b111111010011100100000110, 24'b111111010100001100000001, 24'b111111100110011011101100, 24'b000000000100101011001010, 24'b000000100100000111001000, 24'b000000111000010001110110, 24'b000000110111100010100001, 24'b000000011111000011010110, 24'b111111110100110010001000, 24'b111111000110101010111101, 24'b111110100110111101110100, 24'b111110100110101110000101, 24'b111111010000000110001001, 24'b000000100010010100111110, 24'b000010010000110000001000, 24'b000100000101011001111110, 24'b000101100110100100101110, 24'b000110011101101101110000, 24'b000110011101101101110000, 24'b000101100110100100101110, 24'b000100000101011001111110, 24'b000010010000110000001000, 24'b000000100010010100111110, 24'b111111010000000110001001, 24'b111110100110101110000101, 24'b111110100110111101110100, 24'b111111000110101010111101, 24'b111111110100110010001000, 24'b000000011111000011010110, 24'b000000110111100010100001, 24'b000000111000010001110110, 24'b000000100100000111001000, 24'b000000000100101011001010, 24'b111111100110011011101100, 24'b111111010100001100000001, 24'b111111010011100100000110, 24'b111111100011100010001000, 24'b111111111101010010110111, 24'b000000010111000001111110, 24'b000000100111011110101001, 24'b000000101001000100110101, 24'b000000011011101010000010, 24'b000000000100010000000111, 24'b111111101011001010010100, 24'b111111011001000100000100, 24'b111111010100001001011011, 24'b111111011110001100000000, 24'b111111110100000111100101, 24'b000000001111001000011100, 24'b000000100110110110110100, 24'b000000110011110111101110, 24'b000000110001110001100011, 24'b000000100000001111100100, 24'b000000000010110111000100, 24'b111111011111111001001101, 24'b111110111110011111001000, 24'b111110100100110100101100, 24'b111110010110110010010110, 24'b111110010101011000011000, 24'b111110011110111101100101, 24'b111110110000000100110101, 24'b111111000100100100001011, 24'b111111011000100111111010, 24'b111111101001100000111101, 24'b111111110101110111110011, 24'b111111111101100101100110, 24'b000000000001011100010010, 24'b000000000010101000100000, 24'b000000000010010111000001, 24'b000000000001100011011110, 24'b000000000000110001111111, 24'b000000000000010010001100};


// Pipeline registers for MAC (Multiply-Accumulate) chain
// Each stage holds the running sum of products up to that tap.
reg signed [DATA_OUT_WIDTH-1:0] pipeline [0:TAP_COUNT-1];

integer i, j;


//-----------------------------------------------------------
// Tap Coefficient Initialization
//-----------------------------------------------------------
//initial begin
// $readmemb("lpFilterTapsBinarySigned.txt", taps);
//end

//-----------------------------------------------------------
// Delay Line (Shift Register)
//-----------------------------------------------------------
always @(posedge clk or negedge reset_n) begin
    if (!reset_n) begin
        for (i = 0; i < TAP_COUNT; i = i + 1)
            delay[i] <= 0;
    end else begin
        // Shift the delay line: new sample enters at delay[0]
        for (i = 1; i < TAP_COUNT; i = i + 1)
            delay[i] <= delay[i-1];
        delay[0] <= data_in;
    end
end

//-----------------------------------------------------------
// Pipelined MAC Operation
//-----------------------------------------------------------
// Each stage j adds the product of delay[j] and taps[j] to the running sum.


    
        always @(posedge clk or negedge reset_n) begin
            if (!reset_n) begin
for (j = 0; j < TAP_COUNT; j = j + 1)
                pipeline[j] <= 0;
    end
            else begin
pipeline[0] <=  data_in * taps[0];
for (j = 0; j < TAP_COUNT; j = j + 1)
                pipeline[j+1] <= (delay[j] * taps[j+1]);
    end
        end



//-----------------------------------------------------------
// Final Output Register
//-----------------------------------------------------------

always @(posedge clk or negedge reset_n) begin
    if (!reset_n)
        data_out <= 0;
    else begin
  // Compute filter output
        data_out <= 0;
        for (i = 0; i < TAP_COUNT; i = i + 1) begin
            data_out <= data_out + pipeline[i];
        end
 end
end
endmodule
