module FIR_Filter_L2_Top 
#(
    parameter DATA_IN_WIDTH  = 16,
    parameter DATA_OUT_WIDTH = 64,
    parameter TAP_WIDTH      = 24,
    parameter TAP_COUNT      = 54
)
(
    input wire                               clk,
    input wire                               reset_n,
    input wire   signed [DATA_IN_WIDTH-1:0]  data_in_1,
	 input wire   signed [DATA_IN_WIDTH-1:0]  data_in_2,
    output reg   signed [DATA_OUT_WIDTH-1:0] data_out_1,
	 output reg   signed [DATA_OUT_WIDTH-1:0] data_out_2
);

//input side of diagram
reg [DATA_IN_WIDTH-1:0] data_sum;
assign data_sum = data_in_1 + data_in_2;

// Coefficient values for each tap (to be copied and pasted)
localparam signed [TAP_WIDTH-1:0] H0_taps [0:TAP_COUNT-1] = '{24'b000000000000010010001100, 24'b000000000001100011011110, 24'b000000000010101000100000, 24'b111111111101100101100110, 24'b111111101001100000111101, 24'b111111000100100100001011, 24'b111110011110111101100101, 24'b111110010110110010010110, 24'b111110111110011111001000, 24'b000000000010110111000100, 24'b000000110001110001100011, 24'b000000100110110110110100, 24'b111111110100000111100101, 24'b111111010100001001011011, 24'b111111101011001010010100, 24'b000000011011101010000010, 24'b000000100111011110101001, 24'b111111111101010010110111, 24'b111111010011100100000110, 24'b111111100110011011101100, 24'b000000100100000111001000, 24'b000000110111100010100001, 24'b111111110100110010001000, 24'b111110100110111101110100, 24'b111111010000000110001001, 24'b000010010000110000001000, 24'b000101100110100100101110, 24'b000110011101101101110000, 24'b000100000101011001111110, 24'b000000100010010100111110, 24'b111110100110101110000101, 24'b111111000110101010111101, 24'b000000011111000011010110, 24'b000000111000010001110110, 24'b000000000100101011001010, 24'b111111010100001100000001, 24'b111111100011100010001000, 24'b000000010111000001111110, 24'b000000101001000100110101, 24'b000000000100010000000111, 24'b111111011001000100000100, 24'b111111011110001100000000, 24'b000000001111001000011100, 24'b000000110011110111101110, 24'b000000100000001111100100, 24'b111111011111111001001101, 24'b111110100100110100101100, 24'b111110010101011000011000, 24'b111110110000000100110101, 24'b111111011000100111111010, 24'b111111110101110111110011, 24'b000000000001011100010010, 24'b000000000010010111000001, 24'b000000000000110001111111};

localparam signed [TAP_WIDTH-1:0] H1_taps [0:TAP_COUNT-1] = '{24'b000000000000110001111111, 24'b000000000010010111000001, 24'b000000000001011100010010, 24'b111111110101110111110011, 24'b111111011000100111111010, 24'b111110110000000100110101, 24'b111110010101011000011000, 24'b111110100100110100101100, 24'b111111011111111001001101, 24'b000000100000001111100100, 24'b000000110011110111101110, 24'b000000001111001000011100, 24'b111111011110001100000000, 24'b111111011001000100000100, 24'b000000000100010000000111, 24'b000000101001000100110101, 24'b000000010111000001111110, 24'b111111100011100010001000, 24'b111111010100001100000001, 24'b000000000100101011001010, 24'b000000111000010001110110, 24'b000000011111000011010110, 24'b111111000110101010111101, 24'b111110100110101110000101, 24'b000000100010010100111110, 24'b000100000101011001111110, 24'b000110011101101101110000, 24'b000101100110100100101110, 24'b000010010000110000001000, 24'b111111010000000110001001, 24'b111110100110111101110100, 24'b111111110100110010001000, 24'b000000110111100010100001, 24'b000000100100000111001000, 24'b111111100110011011101100, 24'b111111010011100100000110, 24'b111111111101010010110111, 24'b000000100111011110101001, 24'b000000011011101010000010, 24'b111111101011001010010100, 24'b111111010100001001011011, 24'b111111110100000111100101, 24'b000000100110110110110100, 24'b000000110001110001100011, 24'b000000000010110111000100, 24'b111110111110011111001000, 24'b111110010110110010010110, 24'b111110011110111101100101, 24'b111111000100100100001011, 24'b111111101001100000111101, 24'b111111111101100101100110, 24'b000000000010101000100000, 24'b000000000001100011011110, 24'b000000000000010010001100};

localparam signed [TAP_WIDTH-1:0] H0_H1_taps [0:TAP_COUNT-1] = '{24'b000000000001000100001011, 24'b000000000011111010011111, 24'b000000000100000100110010, 24'b111111110011011101011001, 24'b111111000010001000110111, 24'b111101110100101001000000, 24'b111100110100010101111101, 24'b111100111011100111000010, 24'b111110011110011000010101, 24'b000000100011000110101000, 24'b000001100101101001010001, 24'b000000110101111111010000, 24'b111111010010010011100101, 24'b111110101101001101011111, 24'b111111101111011010011011, 24'b000001000100101110110111, 24'b000000111110100000100111, 24'b111111100000110100111111, 24'b111110100111110000000111, 24'b111111101011000110110110, 24'b000001011100011000111110, 24'b000001010110100101110111, 24'b111110111011011101000101, 24'b111101001101101011111001, 24'b111111110010011011000111, 24'b000110010110001010000110, 24'b001100000100010010011110, 24'b001100000100010010011110, 24'b000110010110001010000110, 24'b111111110010011011000111, 24'b111101001101101011111001, 24'b111110111011011101000101, 24'b000001010110100101110111, 24'b000001011100011000111110, 24'b111111101011000110110110, 24'b111110100111110000000111, 24'b111111100000110100111111, 24'b000000111110100000100111, 24'b000001000100101110110111, 24'b111111101111011010011011, 24'b111110101101001101011111, 24'b111111010010010011100101, 24'b000000110101111111010000, 24'b000001100101101001010001, 24'b000000100011000110101000, 24'b111110011110011000010101, 24'b111100111011100111000010, 24'b111100110100010101111101, 24'b111101110100101001000000, 24'b111111000010001000110111, 24'b111111110011011101011001, 24'b000000000100000100110010, 24'b000000000011111010011111, 24'b000000000001000100001011};




//Data out for sub parallel filters
reg [DATA_OUT_WIDTH-1:0] dataOut_H0;
reg [DATA_OUT_WIDTH-1:0] dataOut_H1;
reg [DATA_OUT_WIDTH-1:0] dataOut_H0H1;

fir_parallel #( .TAPS(H0_taps) ) H0(clk, reset_n, data_in_1, dataOut_H0);
fir_parallel #( .TAPS(H1_taps) ) H1(clk, reset_n, data_in_2, dataOut_H1);
fir_parallel #( .TAPS(H0_H1_taps) ) H0_H1(clk, reset_n, data_sum, dataOut_H0H1);


//output side of diagram:
reg signed [DATA_OUT_WIDTH-1:0] delay;
integer i;
//-----------------------------------------------------------
// Delay Line (for H1)
//-----------------------------------------------------------
always @(posedge clk or negedge reset_n) begin
    if (!reset_n) begin
            delay <= 0;
    end else begin
        // Shift the delay line: new sample enters at delay[0]
        delay <= dataOut_H1;
    end
end


assign data_out_2 = dataOut_H0H1 - dataOut_H1 - dataOut_H0;
assign data_out_1 = dataOut_H0 + delay;

endmodule